--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 

-- ===================================================================

-- coeficientes del filtro y array de muestras (vectores de 9 bits)

-- ===================================================================

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.numeric_std.all;

package filtro_pkg is
	constant Bits_cte_t 	: integer := 24 ; -- agrego 1 bit para tener 23 bits posta  
	constant Bits_x_t		: integer := 8  ;
	constant N_coef		: integer := 21 ; -- el numero de coeficientes del filtro de orden 20

	type x_t is array(integer range <>) of std_logic_vector(Bits_x_t-1 downto 0) ; 
	type cte_t is array(integer range<>) of std_logic_vector(Bits_cte_t-1 downto 0) ; 
	
	-- filtro HAMMING
	constant coefs: cte_t :=  ("000000000000000000000000",                                                       
										"000000001011111111110011",                                                       
										"000000011001111110100111",                                                       
										"000000001111011111101101",                                                       
										"111111001101010000100110",                                                       
										"111101110011011001100000",                                                       
										"111101111101100000001000",                                                       
										"000001101100101011000000",                                                       
										"001000110100101100000000",                                                       
										"010000000101100001010010",                                                       
										"010011001010111110110001",                                                       
										"010000000101100001010010",                                                       
										"001000110100101100000000",                                                       
										"000001101100101011000000",                                                       
										"111101111101100000001000",                                                       
										"111101110011011001100000",                                                       
										"111111001101010000100110",                                                       
										"000000001111011111101101",                                                       
										"000000011001111110100111",                                                       
										"000000001011111111110011",                                                       
										"000000000000000000000000"); 
	
	-- filtro TRIANGULAR
--	constant coefs: cte_t :=  ("000000000000000000000000",                                                       
--										"000000010110011111010011",                                                      
--										"000000101100100111001111",                                                       
--										"000000010110000101101011",                                                       
--										"111111000010101110100110",                                                       
--										"111101101001111001000100",                                                       
--										"111101111111010101000100",                                                       
--										"000001100111000101001000",                                                       
--										"001000010111010110110011",                                                       
--										"001111110100000000001010",                                                       
--										"010100010000110110000001",                                                       
--										"001111110100000000001010",                                                       
--										"001000010111010110110011",                                                       
--										"000001100111000101001000",                                                       
--										"111101111111010101000100",                                                       
--										"111101101001111001000100",                                                       
--										"111111000010101110100110",                                                       
--										"000000010110000101101011",                                                       
--										"000000101100100111001111",                                                       
--										"000000010110011111010011",                                                      
--										"000000000000000000000000");                                                       

                                                                              


 
end filtro_pkg;
                                                                    
                                                      

                                                                              
                                       

                                                                              


					  
      